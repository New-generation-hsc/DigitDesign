-------------------------------
-- Design Unit : datapath 
-- File Name : datapath.vhd

-- Description : 
-- datapath is the combination of different bus and wire
-- it control all port

-- Author : huangshicai
-- mail : 1309508226@qq.com
-- Revision : Version 0.0 2017/12/19
---------------------------------

entity datapath is
	port (
		clock : std_logic;
	);
end datapath;